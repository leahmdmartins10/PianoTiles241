module PianoTilesMaster(CLOCK_50, KEY, SW, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5,
								VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_N, VGA_SYNC_N, //for the VGA adapter
								VGA_R, VGA_G, VGA_B); //for the VGA adapter
								
								input CLOCK_50;
								
								input [8:0] KEY;
								input [9:0] SW;
								output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
								
								output VGA_CLK;
								output VGA_HS;
								output VGA_VS;
								output VGA_BLANK_N;
								output VGA_SYNC_N;
								output [7:0] VGA_R;
								output [7:0] VGA_G;
								output [7:0] VGA_B;
								
								wire resetn;
								wire startn;
								
								assign resetn = SW[0]; // this will need to be changed for when the inputs are sent
								assign startn = KEY[0] | KEY [1] | // this will need to be changed for when the inputs are sent
								
								wire reset_screen_done, drawdone, wait_done,
										reset_screen_go, draw_go, wait_go, edge_go, offset_inc,
										check_input_done,
										correct,
										incorrect,
										correct_done,
										incorrect_input_done,
										color_line_done, check_in_go,
										correct_go,
										incorrect_input_go,
										color_line_go;
							
							wire [5:0] offset;
							
							wire [2:0] line_0, line_1, line_2, line_3, line_4, line_5, line_6;
							
							// vga adpater inputs
							
							wire vga_en;
							wire draw_en, reset_en;
							assign vga_en = draw_vga_en | reset_vga_en | color_line_go | correct_go | incorrect_input_go;
							
							reg [8:0] x;
							wire [8:0] x_draw, x_reset, x_line, x_correct, x_incorrect;
							reg [7:0] y;
							wire [7:0] y_draw, y_reset, y_line, y_correct, y_incorrect;
							
							wire [2:0] color;
							wire [2:0] color_draw, color_reset;
							
							always @(*) begin
								if(reset_screen_go) begin
									x = x_reset;
									y = y_reset;
									color = color_reset;
								end
								else if(draw_go) begin
									x = x_draw;
									y = y_draw;
									color = color_draw;
								end
								else if(color_line_go) begin
									x = x_line;
									y = y_line;
									color = 3'b100;
								end
								else if(correct_go) begin
									x = x_correct;
									y = y_correct;
									color = 3'b111;
								end
								else if(incorrect_input_go) begin
									x = x_incorrect;
									y = y_incorrect;
									color = 3'b100;
								end
								else begin
									x = 1;
									y = 0;
									color = 3'b111;
								end
							end
							
							vga_adapter VGA(.resetn(resetn)
												 .clock(CLOCK_50),
												 .color(color),
												 .x(x),
												 .y(y),
												 .plot(vga_en),
												 .VGA_R(VGA_R),
												 .VGA_G(VGA_G),
												 .VGA_B(VGA_B),
												 .VGA_HS(VGA_HS),
												 .VGA_VS(VGA_VS),
												 .VGA_BLANK_N(VGA_BLANK_N),
												 .VGA_SYNC_N(VGA_SYNC_N),
												 .VGA_CLK(VGA_CLK));
							defparam VGA.RESOLUTION = "320x240";
							defparam VGA.MONOCHROME = "FALSE";
							defparam VGA.BITS_PERCOLOR_CHANNEL = 1;
							defparam VGA.BACKGROUND_IMAGE = "background.mf";
							
							
							wire [5:0] current_state;
							wire [23:0] Q;
							
							all_draw d0(.clock(CLOCK_50),
											.resetn(resetn),
											.startn(startn),
											.draw_go(draw_go),
											.offset([5:0]),
											.line_0(line_0[2:0]),
											.line_1(line_1[2:0]),
											.line_2(line_2[2:0]),
											.line_3(line_3[2:0]),
											.line_4(line_4[2:0]),
											.line_5(line_5[2:0]),
											.line_6(line_6[2:0]),
											.main_state(current_state[5:0]),
											.all_draw_done(drawdone),
											.vga_enable(draw_vga_enable),
											.xOutput(x_draw[8:0]),
											.yOutput(y_draw[7:0]),
											.colorOutput(color_draw[2:0]));
											
							resetScreen reset(.clock(CLOCK_50),
													.reset_screen_go(reset_screen_go),
													.x(x_reset[8:0]),
													.y(y_reset[7:0]),
													.color(color_reset[2:0]),
													.vga_en(reset_vga_en),
													.resetdone(reset_screen_done));
							
							shift	shiftbitch(.shift(edge_go),
												  .clk(CLOCK_50),
												  .resetn(resetn),
												  .startn(startn),
												  .correct_in(correct_done),
												  .current_st(current_state[5:0]),
												  .line_0(line_0[2:0]),
												  .line_1(line_1[2:0]),												  
												  .line_2(line_2[2:0]),
												  .line_3(line_3[2:0]),	
												  .line_4(line_4[2:0]),
												  .line_5(line_5[2:0]),		
												  .line_6(line_6[2:0]));									  
							
							// missing checking input
							
							scoreRegister scoreboard(.clock(CLOCK_50),
															 .resetn(resetn),
															 .startn(startn),
															 .current_state(current_state),
															 .increment(correct_done),
															 .HEX0(HEX0[6:0]),
															 .HEX1(HEX1[6:0]),
															 .HEX2(HEX2[6:0]),
															 .HEX3(HEX3[6:0]),
															 .HEX4(HEX4[6:0]),
															 .HEX5(HEX5[6:0]),
															 .Q(Q[23:0]));
							
							
							
							
							
							
							
							
							
endmodule
